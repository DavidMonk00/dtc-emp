-- emp_project_decl for the VCU118 minimal example design
--
-- Defines constants for the whole project
--


library IEEE;
use IEEE.STD_LOGIC_1164.all;

use work.emp_framework_decl.all;
use work.emp_device_types.all;

-------------------------------------------------------------------------------
package emp_project_decl is

  constant PAYLOAD_REV        : std_logic_vector(31 downto 0) := X"12345678";
  
  -- Number of LHC bunches 
  constant LHC_BUNCH_COUNT    : integer             := 3564;
  -- Latency buffer size
  constant LB_ADDR_WIDTH      : integer             := 10;

  -- Clock setup
  constant CLOCK_COMMON_RATIO : integer             := 24;
  constant CLOCK_RATIO        : integer             := 8;
  constant CLOCK_AUX_RATIO    : clock_ratio_array_t := (2, 4, 6);

  -- Only used by nullalgo
  constant PAYLOAD_LATENCY : integer             := 5;

  -- mgt -> chk -> buf -> fmt -> (algo) -> (fmt) -> buf -> chk -> mgt -> clk -> altclk
  constant REGION_CONF : region_conf_array_t := (
    0  => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    1  => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    2  => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    3  => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    4  => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    5  => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    6  => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    7  => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    8  => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    9  => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    10 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    11 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    12 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    13 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    14 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    15 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    16 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    17 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    18 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    19 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    20 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    21 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    22 => (no_mgt, no_chk, buf   , no_fmt, no_buf, no_chk, no_mgt, -1, -1),
    23 => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    24 => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    25 => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    26 => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    27 => (no_mgt, no_chk, no_buf, no_fmt, buf   , no_chk, no_mgt, -1, -1),
    ---- Cross-chip
    others => kDummyRegion
    );

end emp_project_decl;
-------------------------------------------------------------------------------
